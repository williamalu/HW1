// (~A~B)

module demorgan4
(
 input A,         // Single bit inputs
 input B,
 output nA,       // Output intermediate completed inputs
 output nB,
 output nAandnB   // Single bit output, (~A~B)
);

   wire nA;
   wire nB;
   not Ainv(nA, A); // Top inverter is named Ainv, takes signal A as input and produces signal nA
   not Binv(nB, B);
   and andgate(nAandnB, nA, nB); // AND gate produces nAandnB from nA and nB

endmodule

